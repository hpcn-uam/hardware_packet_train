--/*******************************************************************************
-- *
-- *
-- *  File:
-- *        precise_timestamp.vhd
-- *
-- *
-- *  Module:
-- *        precise_timestamp
-- *
-- *  Author:
-- *        Mario Ruiz
-- *
-- *
-- *  Copyright (C) 2015 - Mario Ruiz and HPCN-UAM High Performance Computing and Networking
-- *
-- *  Licence:
-- *        This file is part of the HPCN-NetFPGA 10G development base package.
-- *
-- *        This file is free code: you can redistribute it and/or modify it under
-- *        the terms of the GNU Lesser General Public License version 2.0 as
-- *        published by the Free Software Foundation.
-- *
-- *        This package is distributed in the hope that it will be useful, but
-- *        WITHOUT ANY WARRANTY; without even the implied warranty of
-- *        MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- *        Lesser General Public License for more details.
-- *
-- *        You should have received a copy of the GNU Lesser General Public
-- *        License along with the NetFPGA source package.  If not, see
-- *        http://www.gnu.org/licenses/.
-- *
-- */

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity precise_timestamp is
    generic (
                 constant width_counter         : integer := 32;
                 constant max_count             : std_logic_vector := x"3B9ACA00";  -- 1.000.000.000 ns
                 constant high_time_pps         : std_logic_vector := x"05F5E100";  -- 100.000.000 ns
                 constant counter_increment     : integer :=10;                     -- 10ns
                 constant max_count_2           : std_logic_vector := x"1DCD6500";  -- 500.000.000 ns 
                 constant fix_point_width       : integer := 3
            );
	port (
			aclk				:	in 	std_logic;
			aresetn			:	in 	std_logic;

			nanosecond		:	out	std_logic_vector(width_counter-1 downto 0);
			second			:	out	std_logic_vector(width_counter-1 downto 0);		
			correction		:	in 	std_logic_vector(width_counter-1 downto 0);

			updatesec			:	in 	std_logic_vector(width_counter-1 downto 0);
			mode				:	in 	std_logic;
			correction_enable 	:	in 	std_logic;

			pps             	:    in   std_logic;
			pps_sync			:	out  std_logic;  
			pps_internal		:	out	std_logic
			
			
		);
end precise_timestamp;

architecture Behavioral of precise_timestamp is

	component counter is
	generic (
        constant width_counter : integer := 32;
        constant max_count : std_logic_vector := x"3B9ACA00"; -- 1.000.000.000 ns
        constant high_time_pps : std_logic_vector := x"05F5E100"; -- 100.000.000 ns
        constant counter_increment : integer :=10 -- 10ns
            ); 
 	port(
		aclk			: 	in 	std_logic;
		aresetn		: 	in 	std_logic;
		timedrift		:	in 	std_logic_vector (1 downto 0);
		pps			:	in	std_logic;
		pps_internal	:	out	std_logic;		
		second 		:	out	std_logic_vector (width_counter-1 downto 0);
		nanosecond	:	out	std_logic_vector (width_counter-1 downto 0);
		mode			:	in	std_logic;
		updatesec		:	in 	std_logic_vector (width_counter-1 downto 0)
		);
	end component;

	

	component tuning is
	generic (
        constant width_counter : integer := 32;
        constant counter_increment : integer :=10 -- 10ns
            );
	port (
			aclk				: 	in 		std_logic;
			aresetn			:	in		std_logic;
			pps				:	in 		std_logic;
			correction		: 	in 		std_logic_vector(width_counter-1 downto 0);
			timedrift			:	out		std_logic_vector(1 downto 0);
			correction_enable	: 	in 		std_logic
		);
	end component;
	
	

	signal 	nsec_counter,sec_counter		: 	std_logic_vector(width_counter-1 downto 0);
	signal	time_corr	                    :	std_logic_vector(width_counter-1 downto 0 );
	signal    time_drift                    : 	std_logic_vector (1 downto 0);   
	signal	pps_out	                    :	std_logic;
	signal	error_calc	               :	std_logic_vector(width_counter-1 downto 0); 
	signal    correction_calc	          :	std_logic_vector(width_counter-1 downto 0);
	signal    pps_ant_ant				: 	std_logic:='0';
	signal    pps_ant					: 	std_logic:='0';


begin


	CONT : counter 
	    generic map (
         		width_counter       => width_counter,
			max_count           => max_count,
			high_time_pps       => high_time_pps,
			counter_increment   => counter_increment
	    )
	    port map(
			aclk			=> aclk,
			aresetn		=> aresetn,
			timedrift		=> time_drift,	
			pps			=> pps_ant_ant,
			pps_internal	=> pps_out,
			second 		=> sec_counter,
			nanosecond	=> nsec_counter,	
			mode			=> mode,
			updatesec		=> updatesec
	);

	TUN : tuning 
	   generic map (
            	width_counter       => width_counter,
            	counter_increment   => counter_increment
	   )
	
	   port map (
			aclk				=> aclk,
			aresetn			=> aresetn,
			pps				=> pps_ant_ant,
			correction		=> correction,
			timedrift			=> time_drift,
			correction_enable	=> correction_enable
		);

	
	


	process (aclk)						-- synchroniser pps
     begin
            if rising_edge(aclk) then
                pps_ant_ant <= pps_ant;
                pps_ant <= pps;
            end if;
    	end process;    
	



	pps_sync 		<= pps_ant_ant;
	pps_internal 	<= pps_out;
	second    	<= sec_counter;
	nanosecond	<= nsec_counter;


--    time_corr <= correction;
--	error_out <= error_calc;
end Behavioral;




